VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vsdmemsoc
  CLASS BLOCK ;
  FOREIGN vsdmemsoc ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 700.000 ;
  PIN CLK
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END CLK
  PIN OUT[0]
    PORT
      LAYER met2 ;
        RECT 54.830 696.000 55.110 700.000 ;
    END
  END OUT[0]
  PIN OUT[1]
    PORT
      LAYER met2 ;
        RECT 164.770 696.000 165.050 700.000 ;
    END
  END OUT[1]
  PIN OUT[2]
    PORT
      LAYER met2 ;
        RECT 274.710 696.000 274.990 700.000 ;
    END
  END OUT[2]
  PIN OUT[3]
    PORT
      LAYER met2 ;
        RECT 384.650 696.000 384.930 700.000 ;
    END
  END OUT[3]
  PIN OUT[4]
    PORT
      LAYER met2 ;
        RECT 494.590 696.000 494.870 700.000 ;
    END
  END OUT[4]
  PIN OUT[5]
    PORT
      LAYER met2 ;
        RECT 604.530 696.000 604.810 700.000 ;
    END
  END OUT[5]
  PIN OUT[6]
    PORT
      LAYER met2 ;
        RECT 714.470 696.000 714.750 700.000 ;
    END
  END OUT[6]
  PIN OUT[7]
    PORT
      LAYER met2 ;
        RECT 824.410 696.000 824.690 700.000 ;
    END
  END OUT[7]
  PIN OUT[8]
    PORT
      LAYER met2 ;
        RECT 934.350 696.000 934.630 700.000 ;
    END
  END OUT[8]
  PIN OUT[9]
    PORT
      LAYER met2 ;
        RECT 1044.290 696.000 1044.570 700.000 ;
    END
  END OUT[9]
  PIN init_addr[0]
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END init_addr[0]
  PIN init_addr[1]
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END init_addr[1]
  PIN init_addr[2]
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END init_addr[2]
  PIN init_addr[3]
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END init_addr[3]
  PIN init_addr[4]
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END init_addr[4]
  PIN init_addr[5]
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END init_addr[5]
  PIN init_addr[6]
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END init_addr[6]
  PIN init_addr[7]
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END init_addr[7]
  PIN init_data[0]
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END init_data[0]
  PIN init_data[10]
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END init_data[10]
  PIN init_data[11]
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END init_data[11]
  PIN init_data[12]
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END init_data[12]
  PIN init_data[13]
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END init_data[13]
  PIN init_data[14]
    PORT
      LAYER met2 ;
        RECT 516.670 0.000 516.950 4.000 ;
    END
  END init_data[14]
  PIN init_data[15]
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END init_data[15]
  PIN init_data[16]
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END init_data[16]
  PIN init_data[17]
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END init_data[17]
  PIN init_data[18]
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END init_data[18]
  PIN init_data[19]
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END init_data[19]
  PIN init_data[1]
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END init_data[1]
  PIN init_data[20]
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END init_data[20]
  PIN init_data[21]
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END init_data[21]
  PIN init_data[22]
    PORT
      LAYER met2 ;
        RECT 781.630 0.000 781.910 4.000 ;
    END
  END init_data[22]
  PIN init_data[23]
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END init_data[23]
  PIN init_data[24]
    PORT
      LAYER met2 ;
        RECT 847.870 0.000 848.150 4.000 ;
    END
  END init_data[24]
  PIN init_data[25]
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END init_data[25]
  PIN init_data[26]
    PORT
      LAYER met2 ;
        RECT 914.110 0.000 914.390 4.000 ;
    END
  END init_data[26]
  PIN init_data[27]
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END init_data[27]
  PIN init_data[28]
    PORT
      LAYER met2 ;
        RECT 980.350 0.000 980.630 4.000 ;
    END
  END init_data[28]
  PIN init_data[29]
    PORT
      LAYER met2 ;
        RECT 1013.470 0.000 1013.750 4.000 ;
    END
  END init_data[29]
  PIN init_data[2]
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END init_data[2]
  PIN init_data[30]
    PORT
      LAYER met2 ;
        RECT 1046.590 0.000 1046.870 4.000 ;
    END
  END init_data[30]
  PIN init_data[31]
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 4.000 ;
    END
  END init_data[31]
  PIN init_data[3]
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END init_data[3]
  PIN init_data[4]
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END init_data[4]
  PIN init_data[5]
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END init_data[5]
  PIN init_data[6]
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END init_data[6]
  PIN init_data[7]
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END init_data[7]
  PIN init_data[8]
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END init_data[8]
  PIN init_data[9]
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END init_data[9]
  PIN init_en
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END init_en
  PIN reset
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END reset
  PIN vccd1
    PORT
      LAYER met5 ;
        RECT 5.280 486.270 1094.580 487.870 ;
    END
    PORT
      LAYER met4 ;
        RECT 1061.340 75.920 1062.940 508.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 639.450 1094.580 641.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 1094.580 334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 1094.580 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 1094.580 28.330 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 503.600 944.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 80.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 504.220 790.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 79.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 503.600 637.040 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 80.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
  END vccd1
  PIN vssd1
    PORT
      LAYER met4 ;
        RECT 1065.020 75.920 1066.620 508.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 642.750 1094.580 644.350 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 489.570 1094.580 491.170 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 1094.580 337.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 1094.580 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 1094.580 31.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 503.600 947.540 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.940 10.640 947.540 80.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 503.600 793.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 79.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 503.600 640.340 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 79.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 688.400 ;
    END
  END vssd1
  PIN _01562_
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 688.400 ;
    END
  END _01562_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1094.340 688.245 ;
      LAYER met1 ;
        RECT 5.520 10.640 1094.340 688.400 ;
      LAYER met2 ;
        RECT 193.360 81.615 1015.490 486.130 ;
      LAYER met3 ;
        RECT 20.310 81.465 1023.380 493.620 ;
      LAYER met4 ;
        RECT 109.100 80.995 174.240 493.620 ;
        RECT 176.640 80.995 177.540 493.620 ;
        RECT 179.940 80.995 327.840 493.620 ;
        RECT 330.240 80.995 331.140 493.620 ;
        RECT 333.540 80.995 481.440 493.620 ;
        RECT 483.840 80.995 484.740 493.620 ;
        RECT 487.140 80.995 1023.380 493.620 ;
  END
END vsdmemsoc
END LIBRARY

